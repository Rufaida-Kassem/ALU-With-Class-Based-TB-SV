`ifndef MONITOR_ALU
`define MONITOR_ALU
`endif
// remaining code to be added here
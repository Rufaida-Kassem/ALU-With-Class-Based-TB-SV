`ifndef MONITOR_ALU
`define MONITOR_ALU
`endif
// remaining, and top-level alu
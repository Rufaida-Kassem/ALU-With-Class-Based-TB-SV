`ifndef MONITOR_ALU
`define MONITOR_ALU
`include "driver.sv"
`include "interface.sv"
`include "transactions.sv"
`include "score_board.sv"
`endif